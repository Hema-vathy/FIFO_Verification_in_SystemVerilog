///////**********PACKAGE OF FILES**********///////
package pkg;
`include "clk_gen.sv"
`include "rst_gen.sv"
`include "tests.sv"
`include "run_test.sv"
endpackage
